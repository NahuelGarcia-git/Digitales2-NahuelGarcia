library verilog;
use verilog.vl_types.all;
entity multiplicador_signo_otro_vlg_vec_tst is
end multiplicador_signo_otro_vlg_vec_tst;
