-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Nov 02 13:22:05 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY I2C IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        soy : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        sda : IN STD_LOGIC := '0';
        ack : OUT STD_LOGIC;
        hab_dir : OUT STD_LOGIC;
        hab_dat : OUT STD_LOGIC
    );
END I2C;

ARCHITECTURE BEHAVIOR OF I2C IS
    TYPE type_fstate IS (Oscioso,Guarda_dir,R_W,A_C_K,Guarda_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,soy,fin_dir,fin_dato,sda)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            ack <= '0';
            hab_dir <= '0';
            hab_dat <= '0';
        ELSE
            ack <= '0';
            hab_dir <= '0';
            hab_dat <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((sda = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((sda = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    ack <= '0';

                    hab_dir <= '0';

                    hab_dat <= '0';
                WHEN Guarda_dir =>
                    IF ((fin_dir = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= R_W;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_dir;
                    END IF;

                    ack <= '0';

                    hab_dir <= '1';

                    hab_dat <= '0';
                WHEN R_W =>
                    reg_fstate <= A_C_K;

                    ack <= '0';

                    hab_dir <= '0';

                    hab_dat <= '0';
                WHEN A_C_K =>
                    reg_fstate <= Guarda_dato;

                    ack <= '1';

                    hab_dir <= '0';

                    hab_dat <= '0';
                WHEN Guarda_dato =>
                    IF ((fin_dato = '0')) THEN
                        reg_fstate <= Guarda_dato;
                    ELSIF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_dato;
                    END IF;

                    ack <= '0';

                    hab_dir <= '0';

                    hab_dat <= '1';
                WHEN OTHERS => 
                    ack <= 'X';
                    hab_dir <= 'X';
                    hab_dat <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
