-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Oct 28 10:39:07 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY State_machine IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z1 : OUT STD_LOGIC;
        z2 : OUT STD_LOGIC;
        z3 : OUT STD_LOGIC;
        z4 : OUT STD_LOGIC
    );
END State_machine;

ARCHITECTURE BEHAVIOR OF State_machine IS
    TYPE type_fstate IS (G,F,E,D,C,B,A);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
            z4 <= '0';
        ELSE
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
            z4 <= '0';
            CASE fstate IS
                WHEN G =>
                    reg_fstate <= A;

                    IF ((x = x)) THEN
                        z4 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN F =>
                    reg_fstate <= C;

                    IF ((x = x)) THEN
                        z4 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN E =>
                    reg_fstate <= F;

                    IF ((x = x)) THEN
                        z4 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN D =>
                    reg_fstate <= A;

                    IF ((x = x)) THEN
                        z4 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z3 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN C =>
                    IF ((x = '0')) THEN
                        reg_fstate <= D;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    IF ((x = '0')) THEN
                        z4 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z3 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z2 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN B =>
                    reg_fstate <= C;

                    IF ((x = x)) THEN
                        z4 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z3 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = x)) THEN
                        z1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN A =>
                    IF ((x = '1')) THEN
                        reg_fstate <= E;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= B;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    IF ((x = '0')) THEN
                        z4 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z4 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z3 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z3 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z2 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z2 <= '0';
                    END IF;

                    IF ((x = '0')) THEN
                        z1 <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z1 <= '0';
                    END IF;
                WHEN OTHERS => 
                    z1 <= 'X';
                    z2 <= 'X';
                    z3 <= 'X';
                    z4 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
