library verilog;
use verilog.vl_types.all;
entity Multiplicador2x2_vlg_vec_tst is
end Multiplicador2x2_vlg_vec_tst;
