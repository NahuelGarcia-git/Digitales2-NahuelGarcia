library verilog;
use verilog.vl_types.all;
entity Inter_Integrated_Circuit_vlg_vec_tst is
end Inter_Integrated_Circuit_vlg_vec_tst;
