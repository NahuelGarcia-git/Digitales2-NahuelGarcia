library verilog;
use verilog.vl_types.all;
entity esquematico_vlg_check_tst is
    port(
        r0              : in     vl_logic;
        r1              : in     vl_logic;
        r2              : in     vl_logic;
        r3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end esquematico_vlg_check_tst;
