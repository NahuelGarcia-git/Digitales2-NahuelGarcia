library verilog;
use verilog.vl_types.all;
entity Multiplicador2x2_vlg_check_tst is
    port(
        P0              : in     vl_logic;
        P1              : in     vl_logic;
        P2              : in     vl_logic;
        P3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Multiplicador2x2_vlg_check_tst;
