library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiplicador_ca2_testbench is
end entity:

architecture comportamiento of multiplicador_ca2_testbench is

component