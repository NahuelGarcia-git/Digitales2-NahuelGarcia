library verilog;
use verilog.vl_types.all;
entity multiplicador_mod_ca2_vlg_vec_tst is
end multiplicador_mod_ca2_vlg_vec_tst;
