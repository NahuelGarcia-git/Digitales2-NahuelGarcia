library verilog;
use verilog.vl_types.all;
entity State_machine_vlg_vec_tst is
end State_machine_vlg_vec_tst;
