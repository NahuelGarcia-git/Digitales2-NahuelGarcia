library verilog;
use verilog.vl_types.all;
entity I2C_vlg_vec_tst is
end I2C_vlg_vec_tst;
