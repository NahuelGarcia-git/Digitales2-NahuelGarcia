library verilog;
use verilog.vl_types.all;
entity Maquina_estado_vlg_vec_tst is
end Maquina_estado_vlg_vec_tst;
